module CRC32 (
	input							Eth_ON,
	input							Clk_125_MHz,
	input				[7:0]		D_In,
	input							En_CRC,

	output			[31:0]	CRC_out
);

reg	[31:0]	Rg_CRC = 32'hff_ff_ff_ff;

//--------------------------------------------------------------------------//
//----------------------- Функция вычисления CRC32. ------------------------//
//--------------------------------------------------------------------------//
function	[31:0]	NextCRC;
	input	[7:0]		D;
	input	[31:0]	C;
	
	reg	[31:0]	NewCRC;

begin
		NewCRC[0]	= C[24]	^ C[30]	^ D[1]	^ D[7];
		NewCRC[1]	= C[25]	^ C[31]	^ D[0]	^ D[6]	^ C[24]	^ C[30]	^ D[1]	^ D[7];
		NewCRC[2]	= C[26]	^ D[5]	^ C[25]	^ C[31]	^ D[0]	^ D[6]	^ C[24]	^ C[30]	^ D[1]	^ D[7];
		NewCRC[3]	= C[27]	^ D[4]	^ C[26]	^ D[5]	^ C[25]	^ C[31]	^ D[0]	^ D[6];
		NewCRC[4]	= C[28]	^ D[3]	^ C[27]	^ D[4]	^ C[26]	^ D[5]	^ C[24]	^ C[30]	^ D[1]	^ D[7];
		NewCRC[5]	= C[29]	^ D[2]	^ C[28]	^ D[3]	^ C[27]	^ D[4]	^ C[25]	^ C[31]	^ D[0]	^ D[6]	^ C[24]	^ C[30]	^ D[1]	^ D[7];
		NewCRC[6]	= C[30]	^ D[1]	^ C[29]	^ D[2]	^ C[28]	^ D[3]	^ C[26]	^ D[5]	^ C[25]	^ C[31]	^ D[0]	^ D[6];
		NewCRC[7]	= C[31]	^ D[0]	^ C[29]	^ D[2]	^ C[27]	^ D[4]	^ C[26]	^ D[5]	^ C[24]	^ D[7];
		NewCRC[8]	= C[0]	^ C[28]	^ D[3]	^ C[27]	^ D[4]	^ C[25]	^ D[6]	^ C[24]	^ D[7];
		NewCRC[9]	= C[1]	^ C[29]	^ D[2]	^ C[28]	^ D[3]	^ C[26]	^ D[5]	^ C[25]	^ D[6];
		NewCRC[10]	= C[2]	^ C[29]	^ D[2]	^ C[27]	^ D[4]	^ C[26]	^ D[5]	^ C[24]	^ D[7];
		NewCRC[11]	= C[3]	^ C[28]	^ D[3]	^ C[27]	^ D[4]	^ C[25]	^ D[6]	^ C[24]	^ D[7];
		NewCRC[12]	= C[4]	^ C[29]	^ D[2]	^ C[28]	^ D[3]	^ C[26]	^ D[5]	^ C[25]	^ D[6]	^ C[24]	^ C[30]	^ D[1]	^ D[7];
		NewCRC[13]	= C[5]	^ C[30]	^ D[1]	^ C[29]	^ D[2]	^ C[27]	^ D[4]	^ C[26]	^ D[5]	^ C[25]	^ C[31]	^ D[0]	^ D[6];
		NewCRC[14]	= C[6]	^ C[31]	^ D[0]	^ C[30]	^ D[1]	^ C[28]	^ D[3]	^ C[27]	^ D[4]	^ C[26]	^ D[5];
		NewCRC[15]	= C[7]	^ C[31]	^ D[0]	^ C[29]	^ D[2]	^ C[28]	^ D[3]	^ C[27]	^ D[4];
		NewCRC[16]	= C[8]	^ C[29]	^ D[2]	^ C[28]	^ D[3]	^ C[24]	^ D[7];
		NewCRC[17]	= C[9]	^ C[30]	^ D[1]	^ C[29]	^ D[2]	^ C[25]	^ D[6];
		NewCRC[18]	= C[10]	^ C[31]	^ D[0]	^ C[30]	^ D[1]	^ C[26]	^ D[5];
		NewCRC[19]	= C[11]	^ C[31]	^ D[0]	^ C[27]	^ D[4];
		NewCRC[20]	= C[12]	^ C[28]	^ D[3];
		NewCRC[21]	= C[13]	^ C[29]	^ D[2];
		NewCRC[22]	= C[14]	^ C[24]	^ D[7];
		NewCRC[23]	= C[15]	^ C[25]	^ D[6]	^ C[24]	^ C[30]	^ D[1]	^ D[7];
		NewCRC[24]	= C[16]	^ C[26]	^ D[5]	^ C[25]	^ C[31]	^ D[0]	^ D[6];
		NewCRC[25]	= C[17]	^ C[27]	^ D[4]	^ C[26]	^ D[5];
		NewCRC[26]	= C[18]	^ C[28]	^ D[3]	^ C[27]	^ D[4]	^ C[24]	^ C[30]	^ D[1]	^ D[7];
		NewCRC[27]	= C[19]	^ C[29]	^ D[2]	^ C[28]	^ D[3]	^ C[25]	^ C[31]	^ D[0]	^ D[6];
		NewCRC[28]	= C[20]	^ C[30]	^ D[1]	^ C[29]	^ D[2]	^ C[26]	^ D[5];
		NewCRC[29]	= C[21]	^ C[31]	^ D[0]	^ C[30]	^ D[1]	^ C[27]	^ D[4];
		NewCRC[30]	= C[22]	^ C[31]	^ D[0]	^ C[28]	^ D[3];
		NewCRC[31]	= C[23]	^ C[29]	^ D[2];
		
		NextCRC	= NewCRC;
	end
endfunction


//--------------------------------------------------------------------------//
//----------------------- Регистр контрольной суммы. -----------------------//
//--------------------------------------------------------------------------//
always @ (posedge Clk_125_MHz)
begin
	if (!Eth_ON)
		Rg_CRC	<=32'hff_ff_ff_ff;
	else if (En_CRC)
		Rg_CRC	<=NextCRC(D_In,Rg_CRC);
end


assign CRC_out	= ~{Rg_CRC[24], Rg_CRC[25], Rg_CRC[26], Rg_CRC[27], Rg_CRC[28], Rg_CRC[29], Rg_CRC[30], Rg_CRC[31],
						 Rg_CRC[16], Rg_CRC[17], Rg_CRC[18], Rg_CRC[19], Rg_CRC[20], Rg_CRC[21], Rg_CRC[22], Rg_CRC[23],
						 Rg_CRC[8],  Rg_CRC[9],  Rg_CRC[10], Rg_CRC[11], Rg_CRC[12], Rg_CRC[13], Rg_CRC[14], Rg_CRC[15],
						 Rg_CRC[0],  Rg_CRC[1],  Rg_CRC[2],  Rg_CRC[3],  Rg_CRC[4],  Rg_CRC[5],  Rg_CRC[6],  Rg_CRC[7]};
        

endmodule
